
module sum_logic (p,g,s) ;

input p,g ;

output s ;

assign s= p ^ g ;

endmodule
